library verilog;
use verilog.vl_types.all;
entity Parallel_Adder_vlg_vec_tst is
end Parallel_Adder_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity The_Or_Circuit_vlg_check_tst is
    port(
        P               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end The_Or_Circuit_vlg_check_tst;

library verilog;
use verilog.vl_types.all;
entity \Three-Chip-Logic-Circuit\ is
    port(
        K               : out    vl_logic;
        B               : in     vl_logic;
        A               : in     vl_logic
    );
end \Three-Chip-Logic-Circuit\;

library verilog;
use verilog.vl_types.all;
entity Boolean_Logic is
    port(
        Z               : out    vl_logic;
        B               : in     vl_logic;
        A               : in     vl_logic;
        C               : in     vl_logic;
        D               : in     vl_logic
    );
end Boolean_Logic;

library verilog;
use verilog.vl_types.all;
entity Boolean_Logic_vlg_vec_tst is
end Boolean_Logic_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity The_Or_Circuit_vlg_vec_tst is
end The_Or_Circuit_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Boolean_Logic_vlg_check_tst is
    port(
        Z               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Boolean_Logic_vlg_check_tst;
